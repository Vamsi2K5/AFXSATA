`include "./design/incl/sata_wrapper_define.svh"