`define ULTRA_GTH