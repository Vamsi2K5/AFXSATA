`define ULTRA_GTY