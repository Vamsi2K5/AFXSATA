`define GTX