/******************************************Copyright@2025**************************************
                                    AdriftXCore  ALL rights reserved
                        https://github.com/AdriftXCore https://gitee.com/adriftxcore
=========================================FILE INFO.============================================
FILE Name       : sata_link_crc.sv
Last Update     : 2025/04/14 22:53:14
Latest Versions : 1.0
========================================AUTHOR INFO.===========================================
Created by      : zhanghx
Create date     : 2025/04/14 22:53:14
Version         : 1.0
Description     : The CRC value is initialized to 0x52325032 as defined in the Serial ATA specification
                    G(X) = X32 + X26 + X23 + X22 + X16 + X12 + X11 + X10 + X8 + X7 + X5 + X4 +X2 +X + 1 
=======================================UPDATE HISTPRY==========================================
Modified by     : 
Modified date   : 
Version         : 
Description     : 
******************************Licensed under the GPL-3.0 License******************************/
module sata_link_crc(
    input  [31:0]   data_in ,//big-endian
    input           crc_init,
    input           crc_en  ,
    output [31:0]   crc_out ,
    input           rst_n   ,
    input           clk      
);
        reg [31:0] lfsr_q;
        reg [31:0] lfsr_c;
        reg [31:0] crc_data_in;
        assign crc_data_in = {data_in[0+:8],data_in[8+:8],data_in[16+:8],data_in[24+:8]};//little-endian
        assign crc_out ={lfsr_q[0+:8],lfsr_q[8+:8],lfsr_q[16+:8],lfsr_q[24+:8]};
        always @(*) begin
                lfsr_c[0] = lfsr_q[0] ^ lfsr_q[6] ^ lfsr_q[9] ^ lfsr_q[10] ^ lfsr_q[12] ^ lfsr_q[16] ^ lfsr_q[24] ^ lfsr_q[25] ^ lfsr_q[26] ^ lfsr_q[28] ^ lfsr_q[29] ^ lfsr_q[30] ^ lfsr_q[31] ^ crc_data_in[0] ^ crc_data_in[6] ^ crc_data_in[9] ^ crc_data_in[10] ^ crc_data_in[12] ^ crc_data_in[16] ^ crc_data_in[24] ^ crc_data_in[25] ^ crc_data_in[26] ^ crc_data_in[28] ^ crc_data_in[29] ^ crc_data_in[30] ^ crc_data_in[31];
                lfsr_c[1] = lfsr_q[0] ^ lfsr_q[1] ^ lfsr_q[6] ^ lfsr_q[7] ^ lfsr_q[9] ^ lfsr_q[11] ^ lfsr_q[12] ^ lfsr_q[13] ^ lfsr_q[16] ^ lfsr_q[17] ^ lfsr_q[24] ^ lfsr_q[27] ^ lfsr_q[28] ^ crc_data_in[0] ^ crc_data_in[1] ^ crc_data_in[6] ^ crc_data_in[7] ^ crc_data_in[9] ^ crc_data_in[11] ^ crc_data_in[12] ^ crc_data_in[13] ^ crc_data_in[16] ^ crc_data_in[17] ^ crc_data_in[24] ^ crc_data_in[27] ^ crc_data_in[28];
                lfsr_c[2] = lfsr_q[0] ^ lfsr_q[1] ^ lfsr_q[2] ^ lfsr_q[6] ^ lfsr_q[7] ^ lfsr_q[8] ^ lfsr_q[9] ^ lfsr_q[13] ^ lfsr_q[14] ^ lfsr_q[16] ^ lfsr_q[17] ^ lfsr_q[18] ^ lfsr_q[24] ^ lfsr_q[26] ^ lfsr_q[30] ^ lfsr_q[31] ^ crc_data_in[0] ^ crc_data_in[1] ^ crc_data_in[2] ^ crc_data_in[6] ^ crc_data_in[7] ^ crc_data_in[8] ^ crc_data_in[9] ^ crc_data_in[13] ^ crc_data_in[14] ^ crc_data_in[16] ^ crc_data_in[17] ^ crc_data_in[18] ^ crc_data_in[24] ^ crc_data_in[26] ^ crc_data_in[30] ^ crc_data_in[31];
                lfsr_c[3] = lfsr_q[1] ^ lfsr_q[2] ^ lfsr_q[3] ^ lfsr_q[7] ^ lfsr_q[8] ^ lfsr_q[9] ^ lfsr_q[10] ^ lfsr_q[14] ^ lfsr_q[15] ^ lfsr_q[17] ^ lfsr_q[18] ^ lfsr_q[19] ^ lfsr_q[25] ^ lfsr_q[27] ^ lfsr_q[31] ^ crc_data_in[1] ^ crc_data_in[2] ^ crc_data_in[3] ^ crc_data_in[7] ^ crc_data_in[8] ^ crc_data_in[9] ^ crc_data_in[10] ^ crc_data_in[14] ^ crc_data_in[15] ^ crc_data_in[17] ^ crc_data_in[18] ^ crc_data_in[19] ^ crc_data_in[25] ^ crc_data_in[27] ^ crc_data_in[31];
                lfsr_c[4] = lfsr_q[0] ^ lfsr_q[2] ^ lfsr_q[3] ^ lfsr_q[4] ^ lfsr_q[6] ^ lfsr_q[8] ^ lfsr_q[11] ^ lfsr_q[12] ^ lfsr_q[15] ^ lfsr_q[18] ^ lfsr_q[19] ^ lfsr_q[20] ^ lfsr_q[24] ^ lfsr_q[25] ^ lfsr_q[29] ^ lfsr_q[30] ^ lfsr_q[31] ^ crc_data_in[0] ^ crc_data_in[2] ^ crc_data_in[3] ^ crc_data_in[4] ^ crc_data_in[6] ^ crc_data_in[8] ^ crc_data_in[11] ^ crc_data_in[12] ^ crc_data_in[15] ^ crc_data_in[18] ^ crc_data_in[19] ^ crc_data_in[20] ^ crc_data_in[24] ^ crc_data_in[25] ^ crc_data_in[29] ^ crc_data_in[30] ^ crc_data_in[31];
                lfsr_c[5] = lfsr_q[0] ^ lfsr_q[1] ^ lfsr_q[3] ^ lfsr_q[4] ^ lfsr_q[5] ^ lfsr_q[6] ^ lfsr_q[7] ^ lfsr_q[10] ^ lfsr_q[13] ^ lfsr_q[19] ^ lfsr_q[20] ^ lfsr_q[21] ^ lfsr_q[24] ^ lfsr_q[28] ^ lfsr_q[29] ^ crc_data_in[0] ^ crc_data_in[1] ^ crc_data_in[3] ^ crc_data_in[4] ^ crc_data_in[5] ^ crc_data_in[6] ^ crc_data_in[7] ^ crc_data_in[10] ^ crc_data_in[13] ^ crc_data_in[19] ^ crc_data_in[20] ^ crc_data_in[21] ^ crc_data_in[24] ^ crc_data_in[28] ^ crc_data_in[29];
                lfsr_c[6] = lfsr_q[1] ^ lfsr_q[2] ^ lfsr_q[4] ^ lfsr_q[5] ^ lfsr_q[6] ^ lfsr_q[7] ^ lfsr_q[8] ^ lfsr_q[11] ^ lfsr_q[14] ^ lfsr_q[20] ^ lfsr_q[21] ^ lfsr_q[22] ^ lfsr_q[25] ^ lfsr_q[29] ^ lfsr_q[30] ^ crc_data_in[1] ^ crc_data_in[2] ^ crc_data_in[4] ^ crc_data_in[5] ^ crc_data_in[6] ^ crc_data_in[7] ^ crc_data_in[8] ^ crc_data_in[11] ^ crc_data_in[14] ^ crc_data_in[20] ^ crc_data_in[21] ^ crc_data_in[22] ^ crc_data_in[25] ^ crc_data_in[29] ^ crc_data_in[30];
                lfsr_c[7] = lfsr_q[0] ^ lfsr_q[2] ^ lfsr_q[3] ^ lfsr_q[5] ^ lfsr_q[7] ^ lfsr_q[8] ^ lfsr_q[10] ^ lfsr_q[15] ^ lfsr_q[16] ^ lfsr_q[21] ^ lfsr_q[22] ^ lfsr_q[23] ^ lfsr_q[24] ^ lfsr_q[25] ^ lfsr_q[28] ^ lfsr_q[29] ^ crc_data_in[0] ^ crc_data_in[2] ^ crc_data_in[3] ^ crc_data_in[5] ^ crc_data_in[7] ^ crc_data_in[8] ^ crc_data_in[10] ^ crc_data_in[15] ^ crc_data_in[16] ^ crc_data_in[21] ^ crc_data_in[22] ^ crc_data_in[23] ^ crc_data_in[24] ^ crc_data_in[25] ^ crc_data_in[28] ^ crc_data_in[29];
                lfsr_c[8] = lfsr_q[0] ^ lfsr_q[1] ^ lfsr_q[3] ^ lfsr_q[4] ^ lfsr_q[8] ^ lfsr_q[10] ^ lfsr_q[11] ^ lfsr_q[12] ^ lfsr_q[17] ^ lfsr_q[22] ^ lfsr_q[23] ^ lfsr_q[28] ^ lfsr_q[31] ^ crc_data_in[0] ^ crc_data_in[1] ^ crc_data_in[3] ^ crc_data_in[4] ^ crc_data_in[8] ^ crc_data_in[10] ^ crc_data_in[11] ^ crc_data_in[12] ^ crc_data_in[17] ^ crc_data_in[22] ^ crc_data_in[23] ^ crc_data_in[28] ^ crc_data_in[31];
                lfsr_c[9] = lfsr_q[1] ^ lfsr_q[2] ^ lfsr_q[4] ^ lfsr_q[5] ^ lfsr_q[9] ^ lfsr_q[11] ^ lfsr_q[12] ^ lfsr_q[13] ^ lfsr_q[18] ^ lfsr_q[23] ^ lfsr_q[24] ^ lfsr_q[29] ^ crc_data_in[1] ^ crc_data_in[2] ^ crc_data_in[4] ^ crc_data_in[5] ^ crc_data_in[9] ^ crc_data_in[11] ^ crc_data_in[12] ^ crc_data_in[13] ^ crc_data_in[18] ^ crc_data_in[23] ^ crc_data_in[24] ^ crc_data_in[29];
                lfsr_c[10] = lfsr_q[0] ^ lfsr_q[2] ^ lfsr_q[3] ^ lfsr_q[5] ^ lfsr_q[9] ^ lfsr_q[13] ^ lfsr_q[14] ^ lfsr_q[16] ^ lfsr_q[19] ^ lfsr_q[26] ^ lfsr_q[28] ^ lfsr_q[29] ^ lfsr_q[31] ^ crc_data_in[0] ^ crc_data_in[2] ^ crc_data_in[3] ^ crc_data_in[5] ^ crc_data_in[9] ^ crc_data_in[13] ^ crc_data_in[14] ^ crc_data_in[16] ^ crc_data_in[19] ^ crc_data_in[26] ^ crc_data_in[28] ^ crc_data_in[29] ^ crc_data_in[31];
                lfsr_c[11] = lfsr_q[0] ^ lfsr_q[1] ^ lfsr_q[3] ^ lfsr_q[4] ^ lfsr_q[9] ^ lfsr_q[12] ^ lfsr_q[14] ^ lfsr_q[15] ^ lfsr_q[16] ^ lfsr_q[17] ^ lfsr_q[20] ^ lfsr_q[24] ^ lfsr_q[25] ^ lfsr_q[26] ^ lfsr_q[27] ^ lfsr_q[28] ^ lfsr_q[31] ^ crc_data_in[0] ^ crc_data_in[1] ^ crc_data_in[3] ^ crc_data_in[4] ^ crc_data_in[9] ^ crc_data_in[12] ^ crc_data_in[14] ^ crc_data_in[15] ^ crc_data_in[16] ^ crc_data_in[17] ^ crc_data_in[20] ^ crc_data_in[24] ^ crc_data_in[25] ^ crc_data_in[26] ^ crc_data_in[27] ^ crc_data_in[28] ^ crc_data_in[31];
                lfsr_c[12] = lfsr_q[0] ^ lfsr_q[1] ^ lfsr_q[2] ^ lfsr_q[4] ^ lfsr_q[5] ^ lfsr_q[6] ^ lfsr_q[9] ^ lfsr_q[12] ^ lfsr_q[13] ^ lfsr_q[15] ^ lfsr_q[17] ^ lfsr_q[18] ^ lfsr_q[21] ^ lfsr_q[24] ^ lfsr_q[27] ^ lfsr_q[30] ^ lfsr_q[31] ^ crc_data_in[0] ^ crc_data_in[1] ^ crc_data_in[2] ^ crc_data_in[4] ^ crc_data_in[5] ^ crc_data_in[6] ^ crc_data_in[9] ^ crc_data_in[12] ^ crc_data_in[13] ^ crc_data_in[15] ^ crc_data_in[17] ^ crc_data_in[18] ^ crc_data_in[21] ^ crc_data_in[24] ^ crc_data_in[27] ^ crc_data_in[30] ^ crc_data_in[31];
                lfsr_c[13] = lfsr_q[1] ^ lfsr_q[2] ^ lfsr_q[3] ^ lfsr_q[5] ^ lfsr_q[6] ^ lfsr_q[7] ^ lfsr_q[10] ^ lfsr_q[13] ^ lfsr_q[14] ^ lfsr_q[16] ^ lfsr_q[18] ^ lfsr_q[19] ^ lfsr_q[22] ^ lfsr_q[25] ^ lfsr_q[28] ^ lfsr_q[31] ^ crc_data_in[1] ^ crc_data_in[2] ^ crc_data_in[3] ^ crc_data_in[5] ^ crc_data_in[6] ^ crc_data_in[7] ^ crc_data_in[10] ^ crc_data_in[13] ^ crc_data_in[14] ^ crc_data_in[16] ^ crc_data_in[18] ^ crc_data_in[19] ^ crc_data_in[22] ^ crc_data_in[25] ^ crc_data_in[28] ^ crc_data_in[31];
                lfsr_c[14] = lfsr_q[2] ^ lfsr_q[3] ^ lfsr_q[4] ^ lfsr_q[6] ^ lfsr_q[7] ^ lfsr_q[8] ^ lfsr_q[11] ^ lfsr_q[14] ^ lfsr_q[15] ^ lfsr_q[17] ^ lfsr_q[19] ^ lfsr_q[20] ^ lfsr_q[23] ^ lfsr_q[26] ^ lfsr_q[29] ^ crc_data_in[2] ^ crc_data_in[3] ^ crc_data_in[4] ^ crc_data_in[6] ^ crc_data_in[7] ^ crc_data_in[8] ^ crc_data_in[11] ^ crc_data_in[14] ^ crc_data_in[15] ^ crc_data_in[17] ^ crc_data_in[19] ^ crc_data_in[20] ^ crc_data_in[23] ^ crc_data_in[26] ^ crc_data_in[29];
                lfsr_c[15] = lfsr_q[3] ^ lfsr_q[4] ^ lfsr_q[5] ^ lfsr_q[7] ^ lfsr_q[8] ^ lfsr_q[9] ^ lfsr_q[12] ^ lfsr_q[15] ^ lfsr_q[16] ^ lfsr_q[18] ^ lfsr_q[20] ^ lfsr_q[21] ^ lfsr_q[24] ^ lfsr_q[27] ^ lfsr_q[30] ^ crc_data_in[3] ^ crc_data_in[4] ^ crc_data_in[5] ^ crc_data_in[7] ^ crc_data_in[8] ^ crc_data_in[9] ^ crc_data_in[12] ^ crc_data_in[15] ^ crc_data_in[16] ^ crc_data_in[18] ^ crc_data_in[20] ^ crc_data_in[21] ^ crc_data_in[24] ^ crc_data_in[27] ^ crc_data_in[30];
                lfsr_c[16] = lfsr_q[0] ^ lfsr_q[4] ^ lfsr_q[5] ^ lfsr_q[8] ^ lfsr_q[12] ^ lfsr_q[13] ^ lfsr_q[17] ^ lfsr_q[19] ^ lfsr_q[21] ^ lfsr_q[22] ^ lfsr_q[24] ^ lfsr_q[26] ^ lfsr_q[29] ^ lfsr_q[30] ^ crc_data_in[0] ^ crc_data_in[4] ^ crc_data_in[5] ^ crc_data_in[8] ^ crc_data_in[12] ^ crc_data_in[13] ^ crc_data_in[17] ^ crc_data_in[19] ^ crc_data_in[21] ^ crc_data_in[22] ^ crc_data_in[24] ^ crc_data_in[26] ^ crc_data_in[29] ^ crc_data_in[30];
                lfsr_c[17] = lfsr_q[1] ^ lfsr_q[5] ^ lfsr_q[6] ^ lfsr_q[9] ^ lfsr_q[13] ^ lfsr_q[14] ^ lfsr_q[18] ^ lfsr_q[20] ^ lfsr_q[22] ^ lfsr_q[23] ^ lfsr_q[25] ^ lfsr_q[27] ^ lfsr_q[30] ^ lfsr_q[31] ^ crc_data_in[1] ^ crc_data_in[5] ^ crc_data_in[6] ^ crc_data_in[9] ^ crc_data_in[13] ^ crc_data_in[14] ^ crc_data_in[18] ^ crc_data_in[20] ^ crc_data_in[22] ^ crc_data_in[23] ^ crc_data_in[25] ^ crc_data_in[27] ^ crc_data_in[30] ^ crc_data_in[31];
                lfsr_c[18] = lfsr_q[2] ^ lfsr_q[6] ^ lfsr_q[7] ^ lfsr_q[10] ^ lfsr_q[14] ^ lfsr_q[15] ^ lfsr_q[19] ^ lfsr_q[21] ^ lfsr_q[23] ^ lfsr_q[24] ^ lfsr_q[26] ^ lfsr_q[28] ^ lfsr_q[31] ^ crc_data_in[2] ^ crc_data_in[6] ^ crc_data_in[7] ^ crc_data_in[10] ^ crc_data_in[14] ^ crc_data_in[15] ^ crc_data_in[19] ^ crc_data_in[21] ^ crc_data_in[23] ^ crc_data_in[24] ^ crc_data_in[26] ^ crc_data_in[28] ^ crc_data_in[31];
                lfsr_c[19] = lfsr_q[3] ^ lfsr_q[7] ^ lfsr_q[8] ^ lfsr_q[11] ^ lfsr_q[15] ^ lfsr_q[16] ^ lfsr_q[20] ^ lfsr_q[22] ^ lfsr_q[24] ^ lfsr_q[25] ^ lfsr_q[27] ^ lfsr_q[29] ^ crc_data_in[3] ^ crc_data_in[7] ^ crc_data_in[8] ^ crc_data_in[11] ^ crc_data_in[15] ^ crc_data_in[16] ^ crc_data_in[20] ^ crc_data_in[22] ^ crc_data_in[24] ^ crc_data_in[25] ^ crc_data_in[27] ^ crc_data_in[29];
                lfsr_c[20] = lfsr_q[4] ^ lfsr_q[8] ^ lfsr_q[9] ^ lfsr_q[12] ^ lfsr_q[16] ^ lfsr_q[17] ^ lfsr_q[21] ^ lfsr_q[23] ^ lfsr_q[25] ^ lfsr_q[26] ^ lfsr_q[28] ^ lfsr_q[30] ^ crc_data_in[4] ^ crc_data_in[8] ^ crc_data_in[9] ^ crc_data_in[12] ^ crc_data_in[16] ^ crc_data_in[17] ^ crc_data_in[21] ^ crc_data_in[23] ^ crc_data_in[25] ^ crc_data_in[26] ^ crc_data_in[28] ^ crc_data_in[30];
                lfsr_c[21] = lfsr_q[5] ^ lfsr_q[9] ^ lfsr_q[10] ^ lfsr_q[13] ^ lfsr_q[17] ^ lfsr_q[18] ^ lfsr_q[22] ^ lfsr_q[24] ^ lfsr_q[26] ^ lfsr_q[27] ^ lfsr_q[29] ^ lfsr_q[31] ^ crc_data_in[5] ^ crc_data_in[9] ^ crc_data_in[10] ^ crc_data_in[13] ^ crc_data_in[17] ^ crc_data_in[18] ^ crc_data_in[22] ^ crc_data_in[24] ^ crc_data_in[26] ^ crc_data_in[27] ^ crc_data_in[29] ^ crc_data_in[31];
                lfsr_c[22] = lfsr_q[0] ^ lfsr_q[9] ^ lfsr_q[11] ^ lfsr_q[12] ^ lfsr_q[14] ^ lfsr_q[16] ^ lfsr_q[18] ^ lfsr_q[19] ^ lfsr_q[23] ^ lfsr_q[24] ^ lfsr_q[26] ^ lfsr_q[27] ^ lfsr_q[29] ^ lfsr_q[31] ^ crc_data_in[0] ^ crc_data_in[9] ^ crc_data_in[11] ^ crc_data_in[12] ^ crc_data_in[14] ^ crc_data_in[16] ^ crc_data_in[18] ^ crc_data_in[19] ^ crc_data_in[23] ^ crc_data_in[24] ^ crc_data_in[26] ^ crc_data_in[27] ^ crc_data_in[29] ^ crc_data_in[31];
                lfsr_c[23] = lfsr_q[0] ^ lfsr_q[1] ^ lfsr_q[6] ^ lfsr_q[9] ^ lfsr_q[13] ^ lfsr_q[15] ^ lfsr_q[16] ^ lfsr_q[17] ^ lfsr_q[19] ^ lfsr_q[20] ^ lfsr_q[26] ^ lfsr_q[27] ^ lfsr_q[29] ^ lfsr_q[31] ^ crc_data_in[0] ^ crc_data_in[1] ^ crc_data_in[6] ^ crc_data_in[9] ^ crc_data_in[13] ^ crc_data_in[15] ^ crc_data_in[16] ^ crc_data_in[17] ^ crc_data_in[19] ^ crc_data_in[20] ^ crc_data_in[26] ^ crc_data_in[27] ^ crc_data_in[29] ^ crc_data_in[31];
                lfsr_c[24] = lfsr_q[1] ^ lfsr_q[2] ^ lfsr_q[7] ^ lfsr_q[10] ^ lfsr_q[14] ^ lfsr_q[16] ^ lfsr_q[17] ^ lfsr_q[18] ^ lfsr_q[20] ^ lfsr_q[21] ^ lfsr_q[27] ^ lfsr_q[28] ^ lfsr_q[30] ^ crc_data_in[1] ^ crc_data_in[2] ^ crc_data_in[7] ^ crc_data_in[10] ^ crc_data_in[14] ^ crc_data_in[16] ^ crc_data_in[17] ^ crc_data_in[18] ^ crc_data_in[20] ^ crc_data_in[21] ^ crc_data_in[27] ^ crc_data_in[28] ^ crc_data_in[30];
                lfsr_c[25] = lfsr_q[2] ^ lfsr_q[3] ^ lfsr_q[8] ^ lfsr_q[11] ^ lfsr_q[15] ^ lfsr_q[17] ^ lfsr_q[18] ^ lfsr_q[19] ^ lfsr_q[21] ^ lfsr_q[22] ^ lfsr_q[28] ^ lfsr_q[29] ^ lfsr_q[31] ^ crc_data_in[2] ^ crc_data_in[3] ^ crc_data_in[8] ^ crc_data_in[11] ^ crc_data_in[15] ^ crc_data_in[17] ^ crc_data_in[18] ^ crc_data_in[19] ^ crc_data_in[21] ^ crc_data_in[22] ^ crc_data_in[28] ^ crc_data_in[29] ^ crc_data_in[31];
                lfsr_c[26] = lfsr_q[0] ^ lfsr_q[3] ^ lfsr_q[4] ^ lfsr_q[6] ^ lfsr_q[10] ^ lfsr_q[18] ^ lfsr_q[19] ^ lfsr_q[20] ^ lfsr_q[22] ^ lfsr_q[23] ^ lfsr_q[24] ^ lfsr_q[25] ^ lfsr_q[26] ^ lfsr_q[28] ^ lfsr_q[31] ^ crc_data_in[0] ^ crc_data_in[3] ^ crc_data_in[4] ^ crc_data_in[6] ^ crc_data_in[10] ^ crc_data_in[18] ^ crc_data_in[19] ^ crc_data_in[20] ^ crc_data_in[22] ^ crc_data_in[23] ^ crc_data_in[24] ^ crc_data_in[25] ^ crc_data_in[26] ^ crc_data_in[28] ^ crc_data_in[31];
                lfsr_c[27] = lfsr_q[1] ^ lfsr_q[4] ^ lfsr_q[5] ^ lfsr_q[7] ^ lfsr_q[11] ^ lfsr_q[19] ^ lfsr_q[20] ^ lfsr_q[21] ^ lfsr_q[23] ^ lfsr_q[24] ^ lfsr_q[25] ^ lfsr_q[26] ^ lfsr_q[27] ^ lfsr_q[29] ^ crc_data_in[1] ^ crc_data_in[4] ^ crc_data_in[5] ^ crc_data_in[7] ^ crc_data_in[11] ^ crc_data_in[19] ^ crc_data_in[20] ^ crc_data_in[21] ^ crc_data_in[23] ^ crc_data_in[24] ^ crc_data_in[25] ^ crc_data_in[26] ^ crc_data_in[27] ^ crc_data_in[29];
                lfsr_c[28] = lfsr_q[2] ^ lfsr_q[5] ^ lfsr_q[6] ^ lfsr_q[8] ^ lfsr_q[12] ^ lfsr_q[20] ^ lfsr_q[21] ^ lfsr_q[22] ^ lfsr_q[24] ^ lfsr_q[25] ^ lfsr_q[26] ^ lfsr_q[27] ^ lfsr_q[28] ^ lfsr_q[30] ^ crc_data_in[2] ^ crc_data_in[5] ^ crc_data_in[6] ^ crc_data_in[8] ^ crc_data_in[12] ^ crc_data_in[20] ^ crc_data_in[21] ^ crc_data_in[22] ^ crc_data_in[24] ^ crc_data_in[25] ^ crc_data_in[26] ^ crc_data_in[27] ^ crc_data_in[28] ^ crc_data_in[30];
                lfsr_c[29] = lfsr_q[3] ^ lfsr_q[6] ^ lfsr_q[7] ^ lfsr_q[9] ^ lfsr_q[13] ^ lfsr_q[21] ^ lfsr_q[22] ^ lfsr_q[23] ^ lfsr_q[25] ^ lfsr_q[26] ^ lfsr_q[27] ^ lfsr_q[28] ^ lfsr_q[29] ^ lfsr_q[31] ^ crc_data_in[3] ^ crc_data_in[6] ^ crc_data_in[7] ^ crc_data_in[9] ^ crc_data_in[13] ^ crc_data_in[21] ^ crc_data_in[22] ^ crc_data_in[23] ^ crc_data_in[25] ^ crc_data_in[26] ^ crc_data_in[27] ^ crc_data_in[28] ^ crc_data_in[29] ^ crc_data_in[31];
                lfsr_c[30] = lfsr_q[4] ^ lfsr_q[7] ^ lfsr_q[8] ^ lfsr_q[10] ^ lfsr_q[14] ^ lfsr_q[22] ^ lfsr_q[23] ^ lfsr_q[24] ^ lfsr_q[26] ^ lfsr_q[27] ^ lfsr_q[28] ^ lfsr_q[29] ^ lfsr_q[30] ^ crc_data_in[4] ^ crc_data_in[7] ^ crc_data_in[8] ^ crc_data_in[10] ^ crc_data_in[14] ^ crc_data_in[22] ^ crc_data_in[23] ^ crc_data_in[24] ^ crc_data_in[26] ^ crc_data_in[27] ^ crc_data_in[28] ^ crc_data_in[29] ^ crc_data_in[30];
                lfsr_c[31] = lfsr_q[5] ^ lfsr_q[8] ^ lfsr_q[9] ^ lfsr_q[11] ^ lfsr_q[15] ^ lfsr_q[23] ^ lfsr_q[24] ^ lfsr_q[25] ^ lfsr_q[27] ^ lfsr_q[28] ^ lfsr_q[29] ^ lfsr_q[30] ^ lfsr_q[31] ^ crc_data_in[5] ^ crc_data_in[8] ^ crc_data_in[9] ^ crc_data_in[11] ^ crc_data_in[15] ^ crc_data_in[23] ^ crc_data_in[24] ^ crc_data_in[25] ^ crc_data_in[27] ^ crc_data_in[28] ^ crc_data_in[29] ^ crc_data_in[30] ^ crc_data_in[31];
        end // always

        always @(posedge clk or negedge rst_n) begin
                if(!rst_n)begin
                    lfsr_q  <= 32'h52325032;
                end
                else if(crc_init)begin
                    lfsr_q  <= 32'h52325032;
                end
                else begin
                    lfsr_q  <= crc_en ? lfsr_c : lfsr_q;
                end
        end // always
endmodule // crc
