`define WAVES